module hello_ModuleA;
    initial begin
        $display("hello");
    end
endmodule
//# sourceMappingURL=hello.sv.map
